** sch_path: /home/leo/Repositories/ihp-sg13g2_leo_ip__ota5t/xschem/ihp-sg13g2_leo_ip__ota5t_tb.sch
**.subckt ihp-sg13g2_leo_ip__ota5t_tb
I0 VDD Ib 10u
C1 Vout GND 1p m=1
x1 Vp Vn Vout VDD VSS Ib ihp-sg13g2_leo_ip__ota5t
V0 VSS GND 0
V2 VDD GND {vdd}
E1 Vp net2 net1 GND 0.5
E2 Vn net2 net1 GND -0.5
Vdm net1 GND ac 1
Vcm net2 GND {vcm}
**** begin user architecture code


.param vdd=1.5
.param vcm=0.75

.control

    save all

    * operating point
    op

    write ihp-sg13g2_leo_ip__ota5t_tb.raw
    set appendwrite

    * run ac simulation
    ac dec 20 1k 100e6

    * measure parameters
    let vout_mag = abs(v(Vout))
    let vout_phase_margin = phase(v(Vout)) * 180/pi + 180
    meas ac A0 find vout_mag at=1k
    meas ac UGF when vout_mag=1 fall=1
    meas ac PM find vout_phase_margin when vout_mag=1

    write ihp-sg13g2_leo_ip__ota5t_tb.raw
.endc




** IHP models
.lib cornerMOSlv.lib mos_tt
.lib cornerMOShv.lib mos_tt
.lib cornerHBT.lib hbt_typ
.lib cornerRES.lib res_typ


**** end user architecture code
**.ends

* expanding   symbol:  ihp-sg13g2_leo_ip__ota5t.sym # of pins=6
** sym_path: /home/leo/Repositories/ihp-sg13g2_leo_ip__ota5t/xschem/ihp-sg13g2_leo_ip__ota5t.sym
** sch_path: /home/leo/Repositories/ihp-sg13g2_leo_ip__ota5t/xschem/ihp-sg13g2_leo_ip__ota5t.sch
.subckt ihp-sg13g2_leo_ip__ota5t Vp Vn Vout VDD VSS Ib
*.ipin Vp
*.ipin Vn
*.opin Vout
*.iopin VDD
*.iopin VSS
*.ipin Ib
XM10 node Ib VSS VSS sg13_lv_nmos w=2u l=1u ng=2 m=1
XM11 Vout net1 VDD VDD sg13_lv_pmos w=2u l=1u ng=2 m=1
XM1 Ib Ib VSS VSS sg13_lv_nmos w=2u l=1u ng=2 m=1
XM2 net1 net1 VDD VDD sg13_lv_pmos w=2u l=1u ng=2 m=1
XM3 Vout Vn node VSS sg13_lv_nmos w=20u l=0.5u ng=4 m=1
XM4 net1 Vp node VSS sg13_lv_nmos w=20u l=0.5u ng=4 m=1
.ends

.GLOBAL GND
.end
